/*-
 * SPDX-License-Identifier: BSD-2-Clause
 *
 * This software was developed by SRI International and the University of
 * Cambridge Computer Laboratory (Department of Computer Science and
 * Technology) under DARPA contract HR0011-18-C-0016 ("ECATS"), as part of the
 * DARPA SSITH research programme.
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in the
 *    documentation and/or other materials provided with the distribution.
 *
 * THIS SOFTWARE IS PROVIDED BY THE AUTHOR AND CONTRIBUTORS ``AS IS'' AND
 * ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 * IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
 * ARE DISCLAIMED.  IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE LIABLE
 * FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 * DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
 * OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
 * HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
 * LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
 * OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
 * SUCH DAMAGE.
 */

/*
 * This file was generated by the parse_counters.py script
 * 2022-08-17 08:23:32.624905
 */

import ISA_Decls::*;

typedef 115 No_Of_Evts;
typedef 39 No_Of_Selected_Evts;

typedef struct {
	Bit#(Report_Width) evt_NO_EV;
	Bit#(Report_Width) evt_REDIRECT;
	Bit#(Report_Width) evt_TRAP;
	Bit#(Report_Width) evt_BRANCH;
	Bit#(Report_Width) evt_JAL;
	Bit#(Report_Width) evt_JALR;
	Bit#(Report_Width) evt_AUIPC;
	Bit#(Report_Width) evt_LOAD;
	Bit#(Report_Width) evt_STORE;
	Bit#(Report_Width) evt_LR;
	Bit#(Report_Width) evt_SC;
	Bit#(Report_Width) evt_AMO;
	Bit#(Report_Width) evt_SERIAL_SHIFT;
	Bit#(Report_Width) evt_INT_MUL_DIV_REM;
	Bit#(Report_Width) evt_FP;
	Bit#(Report_Width) evt_SC_SUCCESS;
	Bit#(Report_Width) evt_LOAD_WAIT;
	Bit#(Report_Width) evt_STORE_WAIT;
	Bit#(Report_Width) evt_FENCE;
	Bit#(Report_Width) evt_F_BUSY_NO_CONSUME;
	Bit#(Report_Width) evt_D_BUSY_NO_CONSUME;
	Bit#(Report_Width) evt_1_BUSY_NO_CONSUME;
	Bit#(Report_Width) evt_2_BUSY_NO_CONSUME;
	Bit#(Report_Width) evt_3_BUSY_NO_CONSUME;
	Bit#(Report_Width) evt_IMPRECISE_SETBOUND;
	Bit#(Report_Width) evt_UNREPRESENTABLE_CAP;
	Bit#(Report_Width) evt_MEM_CAP_LOAD;
	Bit#(Report_Width) evt_MEM_CAP_STORE;
	Bit#(Report_Width) evt_MEM_CAP_LOAD_TAG_SET;
	Bit#(Report_Width) evt_MEM_CAP_STORE_TAG_SET;
	Bit#(Report_Width) evt_INTERRUPT;
} EventsCore deriving (Bits, FShow);

typedef struct {
	Bit#(Report_Width) evt_LD;
	Bit#(Report_Width) evt_LD_MISS;
	Bit#(Report_Width) evt_LD_MISS_LAT;
	Bit#(Report_Width) evt_TLB;
	Bit#(Report_Width) evt_TLB_MISS;
	Bit#(Report_Width) evt_TLB_MISS_LAT;
	Bit#(Report_Width) evt_TLB_FLUSH;
} EventsL1I deriving (Bits, FShow);

typedef struct {
	Bit#(Report_Width) evt_LD;
	Bit#(Report_Width) evt_LD_MISS;
	Bit#(Report_Width) evt_LD_MISS_LAT;
	Bit#(Report_Width) evt_ST;
	Bit#(Report_Width) evt_ST_MISS;
	Bit#(Report_Width) evt_ST_MISS_LAT;
	Bit#(Report_Width) evt_AMO;
	Bit#(Report_Width) evt_AMO_MISS;
	Bit#(Report_Width) evt_AMO_MISS_LAT;
	Bit#(Report_Width) evt_TLB;
	Bit#(Report_Width) evt_TLB_MISS;
	Bit#(Report_Width) evt_TLB_MISS_LAT;
	Bit#(Report_Width) evt_TLB_FLUSH;
	Bit#(Report_Width) evt_EVICT;
} EventsL1D deriving (Bits, FShow);

typedef struct {
	Bit#(Report_Width) evt_WRITE;
	Bit#(Report_Width) evt_WRITE_MISS;
	Bit#(Report_Width) evt_READ;
	Bit#(Report_Width) evt_READ_MISS;
	Bit#(Report_Width) evt_EVICT;
	Bit#(Report_Width) evt_SET_TAG_WRITE;
	Bit#(Report_Width) evt_SET_TAG_READ;
} EventsTGC deriving (Bits, FShow);

typedef struct {
	Bit#(Report_Width) evt_AW_FLIT;
	Bit#(Report_Width) evt_W_FLIT;
	Bit#(Report_Width) evt_W_FLIT_FINAL;
	Bit#(Report_Width) evt_B_FLIT;
	Bit#(Report_Width) evt_AR_FLIT;
	Bit#(Report_Width) evt_R_FLIT;
	Bit#(Report_Width) evt_R_FLIT_FINAL;
} AXI4_Slave_Events deriving (Bits, FShow);

typedef struct {
	Bit#(Report_Width) evt_AW_FLIT;
	Bit#(Report_Width) evt_W_FLIT;
	Bit#(Report_Width) evt_W_FLIT_FINAL;
	Bit#(Report_Width) evt_B_FLIT;
	Bit#(Report_Width) evt_AR_FLIT;
	Bit#(Report_Width) evt_R_FLIT;
	Bit#(Report_Width) evt_R_FLIT_FINAL;
} AXI4_Master_Events deriving (Bits, FShow);

typedef struct {
	Bit#(Report_Width) evt_LD;
	Bit#(Report_Width) evt_LD_MISS;
	Bit#(Report_Width) evt_LD_MISS_LAT;
	Bit#(Report_Width) evt_ST;
	Bit#(Report_Width) evt_ST_MISS;
	Bit#(Report_Width) evt_TLB;
	Bit#(Report_Width) evt_TLB_MISS;
	Bit#(Report_Width) evt_TLB_FLUSH;
	Bit#(Report_Width) evt_EVICT;
} EventsLL deriving (Bits, FShow);

typedef struct {
	Bit#(Report_Width) evt_RENAMED_INST;
	Bit#(Report_Width) evt_WILD_JUMP;
	Bit#(Report_Width) evt_WILD_EXCEPTION;
} EventsTransExe deriving (Bits, FShow);

typedef struct {
	Maybe#(EventsCore) mab_EventsCore;
	Maybe#(EventsL1I) mab_EventsL1I;
	Maybe#(EventsL1D) mab_EventsL1D;
	Maybe#(EventsTGC) mab_EventsTGC;
	Maybe#(AXI4_Slave_Events) mab_AXI4_Slave_Events;
	Maybe#(AXI4_Master_Events) mab_AXI4_Master_Events;
	Maybe#(EventsLL) mab_EventsLL;
	Maybe#(EventsTransExe) mab_EventsTransExe;
} HPMEvents deriving (Bits, FShow);
