import ContinuousMonitoring_IFC :: *;

(*synthesize*)
module mkContinuousMonitoring(ContinuousMonitoring_IFC);
    let axi_mem = interface AxiMem_IFC;
endmodule 